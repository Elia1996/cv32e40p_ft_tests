// Copyright 2020 Politecnico di Torino.


////////////////////////////////////////////////////////////////////////////////
// Engineer:       Elia Ribaldone - s265613@studenti.polito.it                //
//                                                                            //
// Design Name:    config_pkg                                                 //
// Project Name:   cv32e40p Fault tolernat                                    //
// Language:       SystemVerilog                                              //
//                                                                            //
// Description:   Majority voter of 3                                         //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////

`ifndef CONFIG_PKG
    `define CONFIG_PKG
    package config_pkg;
	

    end package
`endif
